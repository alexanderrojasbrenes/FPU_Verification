import uvm_pkg::*;

module top_hvl();
import uvm_pkg::*;
initial begin 
  run_test();	
end
  
endmodule