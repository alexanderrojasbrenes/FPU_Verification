class scoreboard;
  logic [31:0] store [$];
endclass